module send_serial(
    input  logic       clk, rst,
    input  logic [7:0] data_in,
    output logic       data_out,
    input  logic       we,
    output logic       busy
);
endmodule
