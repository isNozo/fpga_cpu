module send_serial(
    input  logic clk, rst,
    output data_out
);
endmodule
